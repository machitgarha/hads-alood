package types is
    type time_array is array(natural) of time;
end package;
